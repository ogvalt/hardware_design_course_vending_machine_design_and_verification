/*
 *	File: if.svh
 *	
 *	Header file with interface description
 *
*/

`ifndef __DUT_IF__
`define __DUT_IF__

interface dut_interface (
							input clk;
							input rst;
						);

endinterface: dut_interface

`endif //__DUT_IF__

